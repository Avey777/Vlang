module main
// import json

// fn test_sqlquery() {
// 	sqldata := sqlquery('1','1000')
// 	// println(sqldata)
// 	// mut jsonstr := json.encode(sqldata) //将[]map[string]string 数据类型 编码为 json 数据类型
// 	// reponse := request(jsonstr)!
// 	// println(reponse)
// }

fn test_request_sqlquery() {

	request_sqlquery()
}